module DataBusBuffer(
    input out_control_logic_data,
    input read,
    input address,
    input enable_read_register,
    input read_register_isr_or_irr,
    input [7:0] control_logic_data,
    input [7:0] interrupt_mask,
    input [7:0] interrupt_request_register,
    input [7:0] in_service_register,
    output reg [7:0] data_bus_out
);

    always @* begin
        if (out_control_logic_data == 1'b1) begin
            data_bus_out = control_logic_data;
        end
        else if (read == 1'b0) begin
            data_bus_out = 8'bz;
        end
        else if (address == 1'b1) begin
            data_bus_out = interrupt_mask;
        end
        else if ((enable_read_register == 1'b1) && (read_register_isr_or_irr == 1'b0)) begin
            data_bus_out = interrupt_request_register;
        end
        else if ((enable_read_register == 1'b1) && (read_register_isr_or_irr == 1'b1)) begin
            data_bus_out = in_service_register;
        end
        else begin
            data_bus_out = 8'bz;
        end
    end

endmodule